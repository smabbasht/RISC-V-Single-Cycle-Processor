module Instruction_Memory #(
    input  [63:0] Inst_address,
    output [31:0] Instruction
);

    

endmodule